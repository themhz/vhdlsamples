LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY diff_synchronous IS
    PORT (
        D : IN STD_LOGIC;
        clock, reset : IN STD_LOGIC;
        Q : OUT STD_LOGIC := '0'
    );
END diff_synchronous;

ARCHITECTURE behavioral OF diff_synchronous IS
BEGIN
    PROCESS (clock, reset)
    BEGIN
        IF falling_edge(clock) THEN
            IF reset = '1' THEN
                Q <= '0';
                ELSE
                Q <= D;
            END IF;
        END IF;
    END PROCESS;
END behavioral;